library verilog;
use verilog.vl_types.all;
entity aud_to_fft_sv_unit is
end aud_to_fft_sv_unit;
